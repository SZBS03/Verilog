module DRAM(
    input wire clk;
    input wire address;
);